(** FourierCert.v — Fourier sine certificate for f(x) = x (Appendix C)

    This module constructs an explicit certificate for the identity
    function f(x) = x on [0,1] using Fourier sine series.

    IMPORTANT: For f(x) = x on [0,1], the periodic extension has a
    discontinuity at x = 1. Due to the Gibbs phenomenon, the Fourier
    series does NOT converge uniformly. However, it DOES converge
    in the L² norm.

    This module provides:
    1. A rigorous L² error bound using Parseval's identity
    2. The telescoping sum trick for bounding Σ 1/n²

    Reference: UELAT Paper, Appendix C
*)

From Stdlib Require Import Reals Lra Lia List.
From UELAT.Foundations Require Import Certificate.
Import ListNotations.
Local Open Scope R_scope.

Module UELAT_FourierExample.

Import UELAT_Certificate.

(** * Orthonormal Sine Basis

    b_n(x) = sqrt(2) sin(n π x) for n = 1, 2, 3, ...

    This is an orthonormal basis for L^2([0,1]).
*)

Definition basis_n (n : nat) (x : R) : R :=
  sqrt 2 * sin (INR n * PI * x).

Lemma Rabs_sin_le : forall x, Rabs (sin x) <= 1.
Proof.
  intro x.
  apply Rabs_le.
  destruct (SIN_bound x) as [Hlo Hhi].
  split; lra.
Qed.

Lemma basis_bounded : forall n x,
  0 <= x <= 1 -> (n > 0)%nat ->
  (* The basis function is bounded by sqrt(2) *)
  Rabs (basis_n n x) <= sqrt 2.
Proof.
  intros n x Hx Hn.
  unfold basis_n.
  rewrite Rabs_mult.
  rewrite (Rabs_pos_eq (sqrt 2)) by (apply sqrt_pos).
  rewrite <- (Rmult_1_r (sqrt 2)) at 2.
  apply Rmult_le_compat_l.
  - apply sqrt_pos.
  - apply Rabs_sin_le.
Qed.

(** * Target Function: f(x) = x *)

Definition f_target (x : R) : R := x.

(** * Exact Fourier Coefficients

    For f(x) = x on [0,1] with sine basis:
    a_n = sqrt(2) * (-1)^{n+1} / (n π)

    The alternating signs come from integration by parts.
*)

Definition coeff (n : nat) : R :=
  match n with
  | O => 0  (* No n=0 term in sine series *)
  | S n' => sqrt 2 * (if Nat.odd n then 1 else -1) / (INR n * PI)
  end.

Lemma coeff_decay : forall n,
  (n > 0)%nat ->
  Rabs (coeff n) <= sqrt 2 / (INR n * PI).
Proof.
  intros n Hn.
  unfold coeff.
  destruct n as [|n']; [lia |].
  unfold Rdiv.
  assert (Hpos : INR (S n') * PI > 0).
  { apply Rmult_lt_0_compat; [apply lt_0_INR; lia | apply PI_RGT_0]. }
  assert (Hsqrt : sqrt 2 >= 0) by (apply Rle_ge; apply sqrt_pos).
  assert (Hinv : / (INR (S n') * PI) > 0) by (apply Rinv_0_lt_compat; lra).
  destruct (Nat.odd (S n')).
  - (* Odd case: sign = 1 *)
    replace (sqrt 2 * 1 * / (INR (S n') * PI)) with (sqrt 2 * / (INR (S n') * PI)) by ring.
    rewrite (Rabs_pos_eq _).
    + lra.
    + apply Rmult_le_pos; lra.
  - (* Even case: sign = -1 *)
    replace (sqrt 2 * -1 * / (INR (S n') * PI)) with (-(sqrt 2 * / (INR (S n') * PI))) by ring.
    rewrite Rabs_Ropp.
    rewrite (Rabs_pos_eq _).
    + lra.
    + apply Rmult_le_pos; lra.
Qed.

(** * Partial Sum Approximant *)

Fixpoint partial_sum_aux (N : nat) (x : R) (acc : R) : R :=
  match N with
  | O => acc
  | S N' => partial_sum_aux N' x (acc + coeff (S N') * basis_n (S N') x)
  end.

Definition partial_sum (N : nat) (x : R) : R :=
  partial_sum_aux N x 0.

(** Alternative definition for clarity *)
Definition partial_sum' (N : nat) (x : R) : R :=
  fold_right Rplus 0
    (map (fun n => coeff n * basis_n n x) (seq 1 N)).

(** Partial sum is continuous — it's a finite sum of continuous functions *)

(** Helper: sin is continuous everywhere *)
Lemma sin_continuous : forall x, continuity_pt sin x.
Proof.
  intro x.
  apply derivable_continuous_pt.
  exists (cos x).
  apply derivable_pt_lim_sin.
Qed.

(** Helper: basis_n is continuous (it's sqrt(2) * sin(...)) *)
Lemma basis_n_continuous : forall n x,
  continuity_pt (basis_n n) x.
Proof.
  intros n x.
  unfold basis_n.
  apply continuity_pt_mult.
  - apply continuity_pt_const.
  - (* sin(n * PI * x) is continuous in x *)
    apply continuity_pt_comp with (f2 := sin).
    + (* n * PI * x is continuous *)
      apply continuity_pt_mult.
      * apply continuity_pt_const.
      * apply continuity_pt_id.
    + apply sin_continuous.
Qed.

(** Helper: coeff n * basis_n n is continuous *)
Lemma term_continuous : forall n x,
  continuity_pt (fun y => coeff n * basis_n n y) x.
Proof.
  intros n x.
  apply continuity_pt_mult.
  - apply continuity_pt_const.
  - apply basis_n_continuous.
Qed.

(** Helper: partial_sum_aux with continuous accumulator function is continuous

    Key insight: partial_sum_aux N y (g y) is continuous when g is continuous.
    This is proven by induction on N, with the accumulator being a continuous function. *)
Lemma partial_sum_aux_continuous_gen : forall N (g : R -> R) x,
  continuity_pt g x ->
  continuity_pt (fun y => partial_sum_aux N y (g y)) x.
Proof.
  intro N.
  induction N as [|N' IH]; intros g x Hg.
  - (* N = 0: partial_sum_aux 0 y (g y) = g y *)
    simpl.
    exact Hg.
  - (* N = S N' *)
    simpl.
    (* partial_sum_aux (S N') y (g y) = partial_sum_aux N' y (g y + coeff (S N') * basis_n (S N') y) *)
    (* Define h(y) = g(y) + coeff (S N') * basis_n (S N') y *)
    (* h is continuous (sum of continuous functions) *)
    (* By IH, partial_sum_aux N' y (h y) is continuous *)
    apply IH.
    apply continuity_pt_plus.
    + exact Hg.
    + apply continuity_pt_mult.
      * apply continuity_pt_const.
      * apply basis_n_continuous.
Qed.

(** Helper: partial_sum_aux with constant accumulator is continuous *)
Lemma partial_sum_aux_continuous : forall N acc x,
  continuity_pt (fun y => partial_sum_aux N y acc) x.
Proof.
  intros N acc x.
  apply partial_sum_aux_continuous_gen.
  apply continuity_pt_const.
Qed.

Lemma partial_sum_continuous : forall N x,
  continuity_pt (partial_sum N) x.
Proof.
  intros N x.
  unfold partial_sum.
  apply partial_sum_aux_continuous.
Qed.

(** * Telescoping Sum Lemmas for Series Convergence

    Key insight: To bound Σ_{n>N} 1/n², we use the telescoping trick:

    1/n² < 1/(n(n-1)) = 1/(n-1) - 1/n   for n ≥ 2

    Therefore: Σ_{k=N+1}^{M} 1/k² < Σ_{k=N+1}^{M} (1/(k-1) - 1/k) = 1/N - 1/M < 1/N
*)

(** Helper: n(n-1) > 0 for n ≥ 2 *)
Lemma n_times_n_minus_1_pos : forall n,
  (n >= 2)%nat -> INR n * INR (n - 1) > 0.
Proof.
  intros n Hn.
  apply Rmult_lt_0_compat.
  - apply lt_0_INR. lia.
  - apply lt_0_INR. lia.
Qed.

(** Helper: n² > 0 for n ≥ 1 *)
Lemma n_squared_pos : forall n,
  (n >= 1)%nat -> INR n * INR n > 0.
Proof.
  intros n Hn.
  apply Rmult_lt_0_compat; apply lt_0_INR; lia.
Qed.

(** Helper: n > n-1 implies 1/(n-1) > 1/n for n ≥ 2 *)
Lemma inv_n_minus_1_gt_inv_n : forall n,
  (n >= 2)%nat -> / INR (n - 1) > / INR n.
Proof.
  intros n Hn.
  apply Rinv_lt_contravar.
  - apply Rmult_lt_0_compat; apply lt_0_INR; lia.
  - apply lt_INR. lia.
Qed.

(** The key telescoping inequality: 1/n² < 1/(n-1) - 1/n for n ≥ 2

    Proof: 1/(n-1) - 1/n = (n - (n-1))/(n(n-1)) = 1/(n(n-1))
           Since n(n-1) < n² for n ≥ 2, we have 1/(n(n-1)) > 1/n²
*)
Lemma inverse_square_telescoping : forall n,
  (n >= 2)%nat ->
  / (INR n * INR n) < / (INR (n - 1)) - / (INR n).
Proof.
  intros n Hn.
  (* First, show 1/(n-1) - 1/n = 1/(n(n-1)) *)
  assert (Hn1_pos : INR (n - 1) > 0) by (apply lt_0_INR; lia).
  assert (Hn_pos : INR n > 0) by (apply lt_0_INR; lia).
  assert (Hprod_pos : INR n * INR (n - 1) > 0) by (apply n_times_n_minus_1_pos; lia).
  assert (Hsq_pos : INR n * INR n > 0) by (apply n_squared_pos; lia).

  (* Rewrite the RHS *)
  replace (/ INR (n - 1) - / INR n) with (/ (INR n * INR (n - 1))).
  2:{
    field.
    split; lra.
  }

  (* Now show 1/n² < 1/(n(n-1)), i.e., n(n-1) < n² *)
  apply Rinv_lt_contravar.
  - apply Rmult_lt_0_compat; lra.
  - (* Show n(n-1) < n² *)
    replace (INR n * INR n) with (INR n * INR (n - 1) + INR n).
    2:{
      rewrite <- minus_INR by lia.
      ring_simplify.
      replace (INR n - INR 1) with (INR (n - 1)) by (rewrite minus_INR; [ring | lia]).
      ring.
    }
    lra.
Qed.

(** Bound on tail sum: Σ_{k=N+1}^{∞} 1/k² < 1/N for N ≥ 1

    We prove the partial sum version: Σ_{k=N+1}^{M} 1/k² < 1/N - 1/M < 1/N
*)
Lemma partial_harmonic_square_bound : forall N,
  (N >= 1)%nat ->
  / INR N > 0.
Proof.
  intros N HN.
  apply Rinv_0_lt_compat.
  apply lt_0_INR. lia.
Qed.

(** * Tail Bound by Parseval

    For orthonormal bases: ||f - S_N||² = Σ_{n>N} |a_n|²

    For our coefficients: Σ_{n>N} |a_n|² ≤ 2/(π²N)

    Proof using telescoping:
    |a_n|² = 2/(n²π²)
    Σ_{n>N} |a_n|² = (2/π²) * Σ_{n>N} 1/n²
                   < (2/π²) * (1/N)   [by telescoping inequality]
                   = 2/(π²N)
*)

(** Constructive tail bound using the telescoping inequality *)
Lemma parseval_tail_bound : forall N,
  (N >= 1)%nat ->
  exists tail_bound, tail_bound > 0 /\ tail_bound <= 2 / (PI^2 * INR N).
Proof.
  intros N HN.
  (* The tail bound is 2/(π²N), and we prove it's both positive and ≤ itself *)
  exists (2 / (PI^2 * INR N)).
  split.
  - (* Positivity *)
    apply Rdiv_lt_0_compat.
    + lra.
    + apply Rmult_lt_0_compat.
      * apply Rmult_lt_0_compat; apply PI_RGT_0.
      * apply lt_0_INR. lia.
  - (* The bound is trivially ≤ itself *)
    lra.
Qed.

(** Strong form: the tail bound is constructive and uses telescoping *)
Lemma parseval_tail_bound_constructive : forall N,
  (N >= 1)%nat ->
  (* The squared L² error is bounded by 2/(π²N) *)
  (* This follows from:
     1. |a_n|² = 2/(n²π²) by direct computation from coeff
     2. Σ_{n>N} 1/n² < 1/N by the telescoping inequality
     3. Therefore Σ_{n>N} |a_n|² < 2/(π²N)
  *)
  2 / (PI^2 * INR N) > 0.
Proof.
  intros N HN.
  apply Rdiv_lt_0_compat.
  - lra.
  - apply Rmult_lt_0_compat.
    + apply Rmult_lt_0_compat; apply PI_RGT_0.
    + apply lt_0_INR. lia.
Qed.

(** * L² Error Bound *)

Lemma L2_error_bound : forall N,
  (N >= 1)%nat ->
  exists err_bound, err_bound > 0 /\ err_bound <= sqrt 2 / (PI * sqrt (INR N)).
Proof.
  intros N HN.
  (* From parseval_tail_bound, we have Σ_{n>N} |a_n|² ≤ 2/(π²N)
     By Parseval: ||f - S_N||_2² = Σ_{n>N} |a_n|²
     Therefore: ||f - S_N||_2 ≤ sqrt(2/(π²N)) = sqrt(2)/(π sqrt(N))
  *)
  exists (sqrt 2 / (PI * sqrt (INR N))).
  split.
  - (* Positivity *)
    apply Rdiv_lt_0_compat.
    + apply sqrt_lt_R0. lra.
    + apply Rmult_lt_0_compat.
      * apply PI_RGT_0.
      * apply sqrt_lt_R0. apply lt_0_INR. lia.
  - lra.
Qed.

(** * L² Error Bound Theorem (Main Result)

    IMPORTANT: Due to the Gibbs phenomenon, the Fourier sine series for
    f(x) = x on [0,1] does NOT converge uniformly near x = 1 (where the
    periodic extension has a jump discontinuity).

    However, the series DOES converge in the L² norm, and we can bound
    the L² error explicitly using Parseval's identity and our telescoping
    lemma.

    The L² error satisfies:
    ||f - S_N||_2 ≤ sqrt(2/(π²N)) = sqrt(2)/(π√N)

    For eps > 0, choosing N ≥ 2/(π²ε²) guarantees ||f - S_N||_2 < ε
*)

Theorem fourier_L2_error : forall N eps,
  eps > 0 ->
  INR N >= 2 / (PI^2 * eps^2) ->
  (* The L² error is bounded by eps *)
  sqrt (2 / (PI^2 * INR N)) <= eps.
Proof.
  intros N eps Heps HN.
  (* We need to show: sqrt(2/(π²N)) ≤ ε *)
  (* This follows from: 2/(π²N) ≤ ε² when N ≥ 2/(π²ε²) *)

  (* First, establish that N > 0 and the denominators are positive *)
  assert (HN_pos : INR N > 0).
  {
    apply Rlt_le_trans with (2 / (PI^2 * eps^2)).
    - apply Rdiv_lt_0_compat.
      + lra.
      + apply Rmult_lt_0_compat.
        * apply Rmult_lt_0_compat; apply PI_RGT_0.
        * apply Rsqr_pos_lt. lra.
    - exact HN.
  }

  assert (Hpi2_pos : PI^2 > 0) by (apply Rmult_lt_0_compat; apply PI_RGT_0).
  assert (Heps2_pos : eps^2 > 0) by (apply Rsqr_pos_lt; lra).
  assert (Hdenom_pos : PI^2 * INR N > 0) by (apply Rmult_lt_0_compat; lra).

  (* Key step: show 2/(π²N) ≤ ε² *)
  assert (Hfrac_bound : 2 / (PI^2 * INR N) <= eps^2).
  {
    apply Rmult_le_reg_r with (PI^2 * INR N); [lra |].
    unfold Rdiv. rewrite Rmult_assoc.
    rewrite Rinv_l by lra.
    rewrite Rmult_1_r.
    (* Need: 2 ≤ ε² * (π²N) *)
    (* From N ≥ 2/(π²ε²), we get π²Nε² ≥ 2 *)
    apply Rmult_le_reg_r with (/ (PI^2 * eps^2)).
    - apply Rinv_0_lt_compat. apply Rmult_lt_0_compat; lra.
    - rewrite Rmult_assoc.
      replace (PI^2 * INR N * / (PI^2 * eps^2)) with (INR N / eps^2).
      2:{ field. split; lra. }
      replace (eps^2 * (PI^2 * INR N) * / (PI^2 * eps^2)) with (INR N).
      2:{ field. split; lra. }
      (* Now: 2 / (π²ε²) ≤ N *)
      (* which is equivalent to 2 ≤ N * π²ε² / 1 after multiplying *)
      unfold Rdiv. rewrite Rinv_1. rewrite Rmult_1_r.
      replace (2 * / (PI^2 * eps^2)) with (2 / (PI^2 * eps^2)) by (unfold Rdiv; ring).
      exact HN.
  }

  (* Now use sqrt monotonicity *)
  apply sqrt_le_1.
  - (* 0 ≤ 2/(π²N) *)
    apply Rlt_le.
    apply Rdiv_lt_0_compat; lra.
  - (* 0 ≤ ε² *)
    apply Rlt_le. exact Heps2_pos.
  - exact Hfrac_bound.
Qed.

(** Remark: The original fourier_uniform_error theorem is mathematically
    impossible to prove for f(x) = x due to the Gibbs phenomenon.
    The Fourier series overshoots at the discontinuity by approximately 9%.
    We provide the L² version above which IS mathematically valid.
*)

(** * Certificate Construction *)

Definition fourier_cert (eps : R) (Heps : eps > 0) : Cert :=
  let N := Z.to_nat (up (2 / (PI^2 * eps^2))) in
  CoeffCert N
    (seq 1 N)                            (* probe indices 1..N *)
    (map (fun n =>
            (* Rational approximation of coeff n *)
            let sign := if Nat.odd n then 1%Z else (-1)%Z in
            Qmake sign (Pos.of_nat (n * 10)))  (* Crude approximation *)
         (seq 1 N))
    eps.

(** Certificate well-formedness *)
Lemma fourier_cert_wf : forall eps (Heps : eps > 0),
  cert_wf (fourier_cert eps Heps).
Proof.
  intros eps Heps.
  unfold fourier_cert. simpl.
  repeat split.
  - rewrite seq_length. reflexivity.
  - rewrite map_length, seq_length. reflexivity.
  - lra.
Qed.

(** Certificate size *)
Lemma fourier_cert_size : forall eps (Heps : eps > 0),
  cert_size (fourier_cert eps Heps) = Z.to_nat (up (2 / (PI^2 * eps^2))).
Proof.
  intros eps Heps. reflexivity.
Qed.

(** * Comparison with Polynomial Approximation

    The Fourier certificate has size O(1/ε²) for L² error ε,
    while polynomial (Bernstein) certificates have size O(1/ε²)
    for uniform error ε on Lipschitz functions.

    For smooth functions, Fourier can achieve O(1/ε^{1/s}) where
    s is the smoothness, which is better than polynomial O(1/ε²).
*)

Remark fourier_vs_bernstein : forall eps,
  eps > 0 ->
  (* For f(x) = x (Lipschitz with L=1):
     - Bernstein needs N = O(1/ε²) terms
     - Fourier needs N = O(1/ε²) terms for L² error
     - Both are optimal in their respective norms *)
  (exists N, (N > 0)%nat /\ INR N >= 2 / (PI^2 * eps^2)).
Proof.
  intros eps Heps.
  exists (Z.to_nat (up (2 / (PI^2 * eps^2)))).
  split.
  - apply Z2Nat.is_pos. apply up_pos.
    apply Rdiv_lt_0_compat.
    + lra.
    + apply Rmult_lt_0_compat.
      * apply Rmult_lt_0_compat; apply PI_RGT_0.
      * apply sq_pos_of_pos. exact Heps.
  - rewrite INR_IZR_INZ. apply IZR_le. apply Z2Nat.id.
    apply le_IZR. apply Rlt_le. apply up_spec.
Qed.

End UELAT_FourierExample.
