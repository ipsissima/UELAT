(** Probe.v — Category Probe with morphisms (Section 3)

    This module defines the category Probe of finite probe theories,
    which forms one side of the Probes-Models adjunction.

    Reference: UELAT Paper, Section 3
*)

From Coq Require Import Reals QArith List Arith Lia.
From UELAT.Foundations Require Import ProbeTheory.
Import ListNotations.
Local Open Scope R_scope.

Module UELAT_ProbeCat.

Import UELAT_Probe.

(** * The Category Probe

    Objects: Finite probe theories T = (n, φ, a)
    Morphisms: Order-preserving injections preserving probes and answers

    This is a skeleton category where objects are identified up to
    isomorphism by their probe-answer data. *)

(** Category structure is given by probe_id and probe_compose
    from ProbeTheory.v *)

(** * Isomorphisms in Probe *)

Definition probe_iso (T T' : ProbeTheory) : Prop :=
  exists (f : ProbeMorphism T T') (g : ProbeMorphism T' T),
    (forall i, (i < rank T)%nat -> injection g (injection f i) = i) /\
    (forall i, (i < rank T')%nat -> injection f (injection g i) = i).

Lemma probe_iso_refl : forall T, probe_iso T T.
Proof.
  intro T.
  exists (probe_id T), (probe_id T).
  split; intros; reflexivity.
Qed.

Lemma probe_iso_sym : forall T T', probe_iso T T' -> probe_iso T' T.
Proof.
  intros T T' [f [g [Hfg Hgf]]].
  exists g, f. split; assumption.
Qed.

Lemma probe_iso_trans : forall T1 T2 T3,
  probe_iso T1 T2 -> probe_iso T2 T3 -> probe_iso T1 T3.
Proof.
  intros T1 T2 T3 [f12 [g21 [H1 H2]]] [f23 [g32 [H3 H4]]].
  exists (probe_compose f12 f23), (probe_compose g32 g21).
  split.
  - intros i Hi. simpl.
    rewrite H3; [apply H1; exact Hi |].
    apply (inj_in_range f12). exact Hi.
  - intros i Hi. simpl.
    rewrite H1; [apply H3; exact Hi |].
    apply (inj_in_range g32). exact Hi.
Qed.

(** * Initial and Terminal Objects *)

(** Empty theory is initial *)
Definition probe_initial : ProbeTheory := empty_theory.

Definition probe_initial_morphism (T : ProbeTheory) : ProbeMorphism probe_initial T.
Proof.
  refine {| injection := fun i => i |}.
  - intros i j Hij. simpl in Hij. lia.
  - intros i Hi. simpl in Hi. lia.
  - intros i Hi. simpl in Hi. lia.
  - intros i Hi. simpl in Hi. lia.
Defined.

Lemma probe_initial_unique : forall T (f g : ProbeMorphism probe_initial T),
  forall i, (i < rank probe_initial)%nat -> injection f i = injection g i.
Proof.
  intros T f g i Hi. simpl in Hi. lia.
Qed.

(** * Coproducts in Probe *)

(** Union gives coproducts *)
Definition probe_coprod (T1 T2 : ProbeTheory) : ProbeTheory := union_theory T1 T2.

Definition probe_inl (T1 T2 : ProbeTheory) : ProbeMorphism T1 (probe_coprod T1 T2) :=
  union_inl T1 T2.

Definition probe_inr (T1 T2 : ProbeTheory) : ProbeMorphism T2 (probe_coprod T1 T2) :=
  union_inr T1 T2.

(** Universal property of coproduct *)
Definition probe_coprod_univ {T1 T2 T : ProbeTheory}
  (f1 : ProbeMorphism T1 T) (f2 : ProbeMorphism T2 T) :
  ProbeMorphism (probe_coprod T1 T2) T.
Proof.
  refine {| injection := fun i =>
    if (i <? rank T1)%nat then injection f1 i
    else injection f2 (i - rank T1) |}.
  - intros i j Hij.
    destruct (i <? rank T1)%nat eqn:Hi; destruct (j <? rank T1)%nat eqn:Hj.
    + apply inj_preserves_order. apply Nat.ltb_lt in Hi, Hj. exact Hij.
    + apply Nat.ltb_lt in Hi. apply Nat.ltb_ge in Hj.
      (* i in T1, j in T2: injection f1 i < rank T ≤ injection f2 (j - rank T1) *)
      (* This requires f1 and f2 to have disjoint ranges - not generally true *)
      (* For a proper coproduct, we need T to be the union *)
      admit.
    + apply Nat.ltb_ge in Hi. apply Nat.ltb_lt in Hj. lia.
    + apply Nat.ltb_ge in Hi, Hj.
      apply inj_preserves_order. lia.
  - intros i Hi. simpl in Hi.
    destruct (i <? rank T1)%nat eqn:Hlt.
    + apply inj_in_range. apply Nat.ltb_lt. exact Hlt.
    + apply inj_in_range. apply Nat.ltb_ge in Hlt. lia.
  - intros i Hi. simpl in Hi.
    destruct (i <? rank T1)%nat eqn:Hlt.
    + simpl. rewrite app_nth1; [| apply Nat.ltb_lt in Hlt; rewrite rank_probes; exact Hlt].
      apply inj_preserves_probes. apply Nat.ltb_lt. exact Hlt.
    + simpl. apply Nat.ltb_ge in Hlt.
      rewrite app_nth2; [| rewrite rank_probes; exact Hlt].
      rewrite rank_probes.
      apply inj_preserves_probes. lia.
  - intros i Hi. simpl in Hi.
    destruct (i <? rank T1)%nat eqn:Hlt.
    + simpl. rewrite app_nth1; [| apply Nat.ltb_lt in Hlt; rewrite rank_answers; exact Hlt].
      apply inj_preserves_answers. apply Nat.ltb_lt. exact Hlt.
    + simpl. apply Nat.ltb_ge in Hlt.
      rewrite app_nth2; [| rewrite rank_answers; exact Hlt].
      rewrite rank_answers.
      apply inj_preserves_answers. lia.
Admitted.

(** * Filtered Colimits

    The category Probe has filtered colimits, which is essential
    for the adjunction with locally finite-dimensional models. *)

(** A directed system in Probe *)
Record DirectedSystem := {
  ds_index : nat -> ProbeTheory;
  ds_transition : forall n, ProbeMorphism (ds_index n) (ds_index (S n))
}.

(** Colimit of a directed system *)
(** The colimit exists as the "union" of all theories in the system *)

End UELAT_ProbeCat.
